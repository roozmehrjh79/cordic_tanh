// FPGA Assignment 4 - Part 1
// Author: Roozmehr Jalilian (97101467)

// CORDIC ROM (Look-up Table)
module cordic_ROM
	#(	// Parameters
		parameter WI = 8,						// fixed-point integer BW
		WF = 16,								// fixed-point fractional BW
		ADDR_DEPTH = 5,							// address depth
		ROM_DEPTH = 1<<ADDR_DEPTH				// ROM depth
	)
	(	// Ports Declaration
		input wire [ADDR_DEPTH-1:0] iAddr,		// input address
		output wire [WI-1:-WF] oQ 				// output (ROM data)
	);

//---------- Wire & Variable Declaration ----------//
		wire [WI-1:-WF] Data [0:ROM_DEPTH-1];	// ROM data
//-------------------------------------------------//

//---------- Continuous Assignments ----------//
		assign Data[0] = 24'h01b78d;
		assign Data[1] = 24'h015aa1;
		assign Data[2] = 24'h00f914;
		assign Data[3] = 24'h008c9f;
		assign Data[4] = 24'h004163;
		assign Data[5] = 24'h00202b;
		assign Data[6] = 24'h001005;
		assign Data[7] = 24'h000801;
		assign Data[8] = 24'h000400;
		assign Data[9] = 24'h000200;
		assign Data[10] = 24'h000100;
		assign Data[11] = 24'h000080;
		assign Data[12] = 24'h000040;
		assign Data[13] = 24'h000020;
		assign Data[14] = 24'h000010;
		assign Data[15] = 24'h000008;
		assign Data[16] = 24'h008000;
		assign Data[17] = 24'h004000;
		assign Data[18] = 24'h002000;
		assign Data[19] = 24'h001000;
		assign Data[20] = 24'h000800;
		assign Data[21] = 24'h000400;
		assign Data[22] = 24'h000200;
		assign Data[23] = 24'h000100;
		assign Data[24] = 24'h000080;
		assign Data[25] = 24'h000040;
		assign Data[26] = 24'h000020;
		assign Data[27] = 24'h000010;
		assign Data[28] = 24'h000008;
		assign Data[29] = 24'h000000;
		assign Data[30] = 24'h000000;
		assign Data[31] = 24'h000000;
		// NOTE: All assignments have been generated by MATLAB code
		
		assign oQ = Data[iAddr];
//--------------------------------------------//

endmodule
